/*`timescale 1ns / 1ps


module aes_tb();

logic CLK = 0;
logic CLR;
logic CK;      //Whenever this is asserted, key is reset
logic [31:0] KEY [7:0];
logic [1:0] KL; 
logic enc_dec;
logic [31:0]state_i[3:0];
logic [31:0]state_o[3:0];
logic CF; 


cipher_unit a(
.CLK(CLK),
.CLR(CLR),
.CK(CK),
.KEY(KEY),
.KL(KL), 
.enc_dec(enc_dec),
.state_i(state_i),
.state_o(state_o),
.CF(CF)
);

always #20 CLK = ~CLK;


// =-=-=-=-=-=-=-=-
logic [31:0] Kzero;     //This is the round key for each round
logic [3:0] round;      //This is the round counter
logic Mux0;             //This controls external input into state
logic Mux1;             //This controls input into BS (byte sub)
logic [1:0]Mux2;        //This controls input into RS(row shift)
logic Mux3;             //This controls input into MC (mix column)
logic Mux4;             //This controls input into ARK (add round key)
logic Mux5;             //This controls input into state (swaps between encryption and decryption flow)
logic Mux6;             //This controls input into ARK (wether MC is skipped or not)
logic [31:0]bso[3:0];
logic [31:0]rso[3:0];
logic [31:0]mco[3:0];
logic [31:0]arko[3:0];
logic [31:0]bsi[3:0];
logic [31:0]rsi[3:0];
logic [31:0]mci[3:0];
logic [31:0]arki[3:0];
logic [3:0]STate;


assign STate = a.s.STATE;
assign Kzero = a.kexp.kout[0];
assign round = a.s.R;
assign Mux0 = a.s.mux0;
assign Mux1 = a.s.mux1;
assign Mux2 = a.s.mux2;
assign Mux3 = a.s.mux3;
assign Mux4 = a.s.mux4;
assign Mux5 = a.s.mux5;
assign Mux6 = a.s.mux6;

assign bsi = a.Bs.state_i;
assign bso = a.Bs.state_o;

assign rsi = a.Rs.state_i;
assign rso = a.Rs.state_o;

assign mci = a.Mc.state_i;
assign mco = a.Mc.state_o;

assign arki = a.Ark.state_i;
assign arko = a.Ark.state_o;


initial 
begin
    //encryption
    enc_dec = 0;//1 is encryption 0 is decryption
    CLR = 1;
    CK = 1;// 1 clears the round keys, 0 does not
    KL = 1;// 0 -> 10 , 1 -> 11 , 2 -> 14

        //USE THIS WHEN TESTING ENCRYPTION, THE NEXT COMMENTED SECTION HAS ITS ENCRYPTED VALUE
  /*  state_i[3] = 32'h2054776F;
    state_i[2] = 32'h4E696E65;
    state_i[1] = 32'h4F6E6520;
    state_i[0] = 32'h54776F20;*/
    /**/
    
    /*  //USE THIS WHEN TESTING DECRYPTION, THE PREVIOUS COMMENTED SECTION HAS ITS DECRYPTED VALUE
    state_i[3] = 32'h1a02d73a;
    state_i[2] = 32'h402299b3;
    state_i[1] = 32'h571420f6;
    state_i[0] = 32'h29c3505f;
    */

/*    
    state_i[0] = 32'hB521EC42;
    state_i[1] = 32'h512227E7;
    state_i[2] = 32'h4B56EFF0;
    state_i[3] = 32'h3A398851;
    
   
    KEY[0] =32'h54686174;
    KEY[1] =32'h73206D79;
    KEY[2] =32'h204B756E;
    KEY[3] =32'h67204675;
    KEY[4] =32'h00000000;
    KEY[5] =32'h00000000;
    KEY[6] =32'h00000000;
    KEY[7] =32'h00000000;
  
    #40

    CLR = 0;
    CK = 0;
    
    #440//          checking stall
    
    #440//          checking encryption
    #40
    #40
    #40
    
    #100



$stop;
$finish;
end



endmodule
*/



`timescale 1ns / 1ps

module aes_tb();

    // Clock and control signals
    logic CLK = 0;
    logic CLR;
    logic CK;      // Key reset
    logic [31:0] KEY [7:0];
    logic [1:0] KL; 
    logic enc_dec;
    logic [31:0] state_i[3:0];
    logic [31:0] state_o[3:0];
    logic CF;

    // Instantiate AES module
    cipher_unit a(
        .CLK(CLK),
        .CLR(CLR),
        .CK(CK),
        .KEY(KEY),
        .KL(KL), 
        .enc_dec(enc_dec),
        .state_i(state_i),
        .state_o(state_o),
        .CF(CF)
    );

    // Clock generation
    always #20 CLK = ~CLK;

    // File handling
    integer infile, outfile;
    integer scanned;
    logic [31:0] word0, word1, word2, word3;
    logic [31:0] plain_i[3:0];
    logic [31:0] cipher_out[3:0];
    logic [31:0] decrypt_out[3:0];

    initial begin
        // ----------------------------
        // Load plaintext and key
        // ----------------------------
        // Example plaintext
        plain_i[3] = 32'h2054776F;
        plain_i[2] = 32'h4E696E65;
        plain_i[1] = 32'h4F6E6520;
        plain_i[0] = 32'h54776F20;

        // AES 256-bit key
        KEY[0] = 32'h54686174;
        KEY[1] = 32'h73206D79;
        KEY[2] = 32'h204B756E;
        KEY[3] = 32'h67204675;
        KEY[4] = 32'h00000000;
        KEY[5] = 32'h00000000;
        KEY[6] = 32'h00000000;
        KEY[7] = 32'h00000000;

        // ----------------------------
        // 1. ENCRYPTION
        // ----------------------------
        enc_dec = 1; // 1 = encryption
        CLR = 1;
        CK = 1;
        KL = 1;      // Key length setting

        #40
        CLR = 0;
        CK = 0;
        #40

        // Apply plaintext to input
        state_i = plain_i;

        // Wait for encryption to complete (CF flag)
        while (CF !== 1) @(posedge CLK);
        @(posedge CLK);

        // Store ciphertext
        cipher_out = state_o;

        $display("Plaintext : %h %h %h %h", plain_i[3], plain_i[2], plain_i[1], plain_i[0]);
        $display("Ciphertext: %h %h %h %h", cipher_out[3], cipher_out[2], cipher_out[1], cipher_out[0]);

        // ----------------------------
        // 2. DECRYPTION
        // ----------------------------
        enc_dec = 0; // 0 = decryption
        state_i = cipher_out;

        // Wait for decryption to complete
        while (CF !== 1) @(posedge CLK);
        @(posedge CLK);

        decrypt_out = state_o;

        $display("Decrypted : %h %h %h %h", decrypt_out[3], decrypt_out[2], decrypt_out[1], decrypt_out[0]);

        // ----------------------------
        // 3. CHECK RESULT
        // ----------------------------
        if (decrypt_out === plain_i)
            $display("SUCCESS: Decrypted output matches original plaintext!");
        else
            $display("ERROR: Decrypted output does NOT match plaintext!");

        #100 $stop;
        $finish;
    end

endmodule














